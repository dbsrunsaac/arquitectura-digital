library ieee;
use ieee.std_logid_1164.all;

entity memory_ram is
port(
	
);
end entity;


architecture Arch of memory_ram is 
begin
	
	
end architecture;