-- Librerías
library ieee;
use ieee.std_logic_1164.all;

entity rom256x8 is
port(
	address : in std_logic_vector(7 downto 0);
	en : in std_logic;
	
);
end entity;

architecture arch of rom256x8 is

begin
	
end;
